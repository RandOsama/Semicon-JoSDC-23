/*module Inst_mem(addr,Inst26_31,Inst21_25,Inst16_20,Inst11_15,Inst0_15,Inst0_5,Inst0_25);

	input [31:0] addr;
	
	output[15:0] Inst0_15;
	output [4:0] Inst11_15,Inst16_20,Inst21_25;
	output [5:0] Inst26_31 , Inst0_5;
	output [25:0] Inst0_25;
	
	reg [31:0] memory [1023:0];
	
	reg [31:0] out;
	
	always@(addr)
		out = memory[addr];
		
	assign Inst0_15 = out[15:0];
	assign Inst11_15 = out[15:11];
	assign Inst16_20 = out[20:16];
	assign Inst21_25 = out[25:21];
	assign Inst26_31 = out[31:26];
	assign Inst0_25 = out[25:0];
	assign Inst0_5 = out[5:0];
	
endmodule*/


module Inst_mem(addr,Inst);

	input [31:0] addr;
	output [31:0]Inst;
	
	reg [31:0] mem [1023:0];
	
	initial begin
	/*
		// arrays1
			mem[0]=32'b10001100000010000000000000000000;
			mem[1]=32'b10001100000010010000000000001000;
			mem[2]=32'b10001100000010100000000000010100;
			mem[3]=32'b10001100000010110000000000000010;
	*/
	/*
		// arrays2
			mem[0]=32'b10001100000000010000000000000010;
			mem[1]=32'b00000000000000010000100010000000;
			mem[2]=32'b10101100000000010000000000000001;
			mem[3]=32'b10001100000000100000000000000001;
			mem[4]=32'b10001100000000110000000000000100;
			mem[5]=32'b00000000000000110001100001000000;
			mem[6]=32'b10101100000000110000000000000011;
			mem[7]=32'b10001100000001000000000000000011;
	*/
	/*
		// Arithmetic Operations
			mem[0]=32'b10001111100010000000000000000000;
			mem[1]=32'b10001111100010010000000000000001;
			mem[2]=32'b00000001000010010100000000100000;
			mem[3]=32'b10001111100010100000000000000010;
			mem[4]=32'b00000001010010100101000000100000;
			mem[5]=32'b00000001000010100100000000100010;
			mem[6]=32'b00100001000010000000000000000001;
			mem[7]=32'b00000000000010000100000000100010;
			
	*/
	/*
		// Conditional statements#1
			mem[0]=32'b00000001000000000100000000100000;
			mem[1]=32'b00100001001010010000000000010000;
			mem[2]=32'b00000001000010010101000000100010;
			mem[3]=32'b00000000000010100101100000101010;
			
			mem[4]=32'b00100000000011000000000000000001;
			mem[5]=32'b00010001100010110000000000000010;
			mem[6]=32'b00100001000010000000000000000001;
			mem[7]=32'b00001000000000000000000000000010;
			mem[8]=32'b00000001001000000110100000100000;
			mem[9]=32'b00100000000011100000000000011011;
			mem[10]=32'b00110001110011100000000000010111;
	*/
	/*	
		// Conditional statements#1
			//case a = 2
				//mem[0]=32'b00100000000000010000000000000010;
			//case a = 6
				mem[0]=32'b00100000000000010000000000000110;
			mem[1]=32'b00100000000000100000000000000010;
			mem[2]=32'b00100000010000110000000000000011;
			mem[3]=32'b00000000001000110010000000101010;
			mem[4]=32'b00010000000001000000000000000010;
			mem[5]=32'b00100000001000010000000000000001;
			mem[6]=32'b00001000000000000000000000001000;
			mem[7]=32'b00100000001000010000000000000010;
			mem[8]=32'b00000000010000010001000000100000;
	*/
		
		// while Loop
			mem[0]=32'b00000000000000000000100000100000;
			mem[1]=32'b00000000000000000001000000100000;
			mem[2]=32'b00100000000010010000000001100100;
			mem[3]=32'b00010001001000010000000000000010;
			mem[4]=32'b00100000001000010000000000000001;
			mem[5]=32'b00001000000000000000000000000011;
			mem[6]=32'b00000000000000000001100000100000;
			mem[7]=32'b00010000000000001111111111111111;

		
	end
	
	assign Inst = mem[addr];
	//initial 
	//begin 
	//$readmemh("C:/Users/Rand5/OneDrive/Desktop/Rand/JOSDC_23/final/instructions.txt",mem);	
	//end 
endmodule 